module shift_reg_tb ;
  reg clk ; 
  reg clr ;
  reg dir ;  
  reg [ N-1 : 0 ] q;
