`timescale 1ns / 1ps 

module uart_tb () ; 

`include " uart_tx.v"
`include " uart_rx.v"

  

  
  
