module shift_reg_tb (
