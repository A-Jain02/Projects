`timescale 1ns / 1ps

module TC_calculator ; 

  
  
