`timescale 1ns / 1ps

module TC_calculator ; 
  reg [3:0] a ;
  reg [3:0] b ;  
  reg [2:0] oper ; 

  wire [7:0] out; 
  

  
  
