`timescale 10ns/10ps



module True_DPR ( clk , en_a , en_b ,
