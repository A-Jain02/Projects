module shift_reg_tb ;
  reg [ N-1 : 0 ] a;
  reg [ 
