`timescale 1ns / 1ps

module uart_rx #(
